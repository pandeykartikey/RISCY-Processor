`timescale 1ns / 1ps

module InstructionMemoryModule(
    input wire clk,
    input wire [31:0] instructionAddress,
    output wire [31:0] instruction
    );


endmodule